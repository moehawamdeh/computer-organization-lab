package constants is
	constant BUS_WIDTH : integer := 8;
end constants;
